// -----------------------------------------------------------------------------
// 文件名: params.vh
// 描述: 定义加速器的全局参数
// -----------------------------------------------------------------------------

`ifndef PARAMS_VH
`define PARAMS_VH

// -----------------------------------------------------------------------------
// 阵列维度定义 (物理维度)
// -----------------------------------------------------------------------------
// 为了适应 Zynq-7020 的 DSP资源 (220个)，我们选择 12x16
// 注意：宏定义不加分号
`define ARRAY_ROW 12
`define ARRAY_COL 16

// -----------------------------------------------------------------------------
// 数据位宽定义
// -----------------------------------------------------------------------------
`define DATA_WIDTH    8
`define ACC_WIDTH     32
`define AXI_DATA_WIDTH 64

// -----------------------------------------------------------------------------
// 默认计数器阈值 (可运行时配置)
// -----------------------------------------------------------------------------
// DeiT-Tiny Hidden Dimension = 192.
// 我们假设每次计算处理一个 Tile 的 K 维度。
`define DEFAULT_K_DIM 192 

`endif