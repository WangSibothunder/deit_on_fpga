// 
`timescale 1ns / 1ps
`include "params.vh"

module deit_core_verify_tb;

    // --- Parameters ---
    parameter CLK_PERIOD = 10.0;
    parameter LATENCY_CFG = 28;
    
    // --- Signals ---
    reg clk, rst_n;
    reg ap_start;
    reg [31:0] cfg_seq_len;
    reg cfg_acc_mode;
    wire ap_done, ap_idle;

    // Buffer Control Signals (From Core)
    wire ctrl_weight_dma_req;   // [CHECK THIS]
    wire ctrl_weight_load_en;   // [CHECK THIS]
    wire ctrl_input_stream_en;

    // Data Interfaces (Simulating AXI Stream)
    reg  [63:0] s_axis_w_tdata;
    reg         s_axis_w_tvalid;
    wire        s_axis_w_tready; // Ignored

    reg  [63:0] s_axis_in_tdata;
    reg         s_axis_in_tvalid;
    
    // Interconnects
    wire [`ARRAY_COL*8-1:0] wbuf_to_core;
    wire [`ARRAY_ROW*8-1:0] ibuf_to_core;
    wire [`ARRAY_COL*32-1:0] out_acc_vec;

    // --- DUT Instantiation ---
    
    // 1. Weight Buffer (Real Module)
    weight_buffer_ctrl u_wbuf (
        .clk(clk), .rst_n(rst_n),
        .s_axis_tdata(s_axis_w_tdata),
        .s_axis_tvalid(s_axis_w_tvalid), // Driven by TB based on DMA Req
        .i_weight_load_en(ctrl_weight_load_en), // Driven by Core (Phase 2)
        .o_weight_vec(wbuf_to_core),
        .i_bank_swap(1'b0)
    );

    // 2. Input Buffer (Real Module)
    input_buffer_ctrl u_ibuf (
        .clk(clk), .rst_n(rst_n),
        .s_axis_tdata(s_axis_in_tdata),
        .s_axis_tvalid(s_axis_in_tvalid),
        .i_rd_en(ctrl_input_stream_en),
        .o_array_vec(ibuf_to_core),
        .i_bank_swap(1'b0)
    );

    // 3. DeiT Core (DUT)
    deit_core #(
        .LATENCY_CFG(LATENCY_CFG),
        .ADDR_WIDTH(8)
    ) u_core (
        .clk(clk), .rst_n(rst_n),
        .ap_start(ap_start),
        .cfg_compute_cycles(cfg_seq_len),
        .cfg_acc_mode(cfg_acc_mode),
        .ap_done(ap_done),
        .ap_idle(ap_idle),
        .in_act_vec(ibuf_to_core),
        .in_weight_vec(wbuf_to_core),
        .out_acc_vec(out_acc_vec),
        .ctrl_weight_dma_req(ctrl_weight_dma_req), // Monitor this!
        .ctrl_weight_load_en(ctrl_weight_load_en), // Monitor this!
        .ctrl_input_stream_en(ctrl_input_stream_en)
    );

    // --- Test Logic ---
    reg [127:0] weight_mem [0:11]; // 12 rows
    reg [95:0]  input_mem  [0:31]; // 32 inputs
    reg [31:0]  load_idx;

    initial begin
        // Init
        clk = 0; rst_n = 0;
        ap_start = 0; cfg_seq_len = 32; cfg_acc_mode = 0;
        s_axis_w_tvalid = 0; s_axis_in_tvalid = 0;
        
        $readmemh("src/test_data_core/weights.mem", weight_mem);
        // Note: Input mem loading skipped for brevity, generated by python
        
        // Reset
        #100 rst_n = 1;
        #20  ap_start = 1; 
        #10  ap_start = 0;

        // [CKPT 1] State: IDLE -> LOAD_W
        wait(ctrl_weight_dma_req == 1);
        $display("[CKPT 1] Phase 1 Started: DMA Req asserted. Time: %t", $time);

        // Feed Weights (Simulate DMA)
        // Need to send 12 rows * 2 beats = 24 beats
        load_idx = 0;
        while (ctrl_weight_dma_req) begin
            @(posedge clk);
            s_axis_w_tvalid = 1;
            // Mock Data: split 128-bit into two 64-bit
            // Simplified: Just sending constant for checking flow
            s_axis_w_tdata = 64'hDEADBEEFCAFEBABE; 
        end
        s_axis_w_tvalid = 0;
        $display("[CKPT 2] Phase 1 Ended: DMA Req deasserted. Time: %t", $time);

        // [CKPT 3] Phase 2: Array Load
        wait(ctrl_weight_load_en == 1);
        $display("[CKPT 3] Phase 2 Started: Array Load asserted. Time: %t", $time);
        
        // Wait for Compute
        wait(ctrl_input_stream_en == 1);
        $display("[CKPT 4] Compute Started. Time: %t", $time);

        wait(ap_done);
        $display("[CKPT 5] DONE Signal Received. Test PASSED. Time: %t", $time);
        $finish;
    end
    
    always #5 clk = ~clk;

endmodule